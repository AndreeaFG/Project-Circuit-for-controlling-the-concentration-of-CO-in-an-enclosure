** Profile: "SCHEMATIC1-param_cc"  [ C:\USERS\SEPTIMIU\DOCUMENTS\DIDACTIC\TCRME\2023\ProiectTCAD-PSpiceFiles\SCHEMATIC1\param_cc.sim ] 

** Creating circuit file "param_cc.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Septimiu\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM Rp 45k 90k 5k 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
